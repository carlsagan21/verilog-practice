// Verilog model of circuit of Figure 3.35 in Digital Systems 5th ed.

module main(A, B, C, D, E);
  parameter WIDTH = 8;

  output D, E;
  input A, B, C;

  wire w1;

  integer i, j;
  integer data[7:0];

endmodule
